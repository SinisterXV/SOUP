library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity digitLUT is
  Port (A: in  std_logic_vector(5 downto 0);
        B: in  std_logic_vector(2 downto 0);
        q: out std_logic_vector(2 downto 0));
end entity;

architecture BEHAVIORAL of digitLUT is
  type LUTtype is array(0 to 511) of std_logic_vector(2 downto 0);

  constant LUT: LUTType := ("000", "000", "001", "001", "001", "001", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "111", "111", "111", "111", "000", "000", 
                            "000", "000", "001", "001", "001", "001", "001", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "111", "111", "111", "111", "111", "000", "000", 
                            "000", "000", "001", "001", "001", "001", "001", "001", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "111", "111", "111", "111", "111", "111", "000", "000", 
                            "000", "000", "001", "001", "001", "001", "001", "001", 
                            "001", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "111", 
                            "111", "111", "111", "111", "111", "111", "000", "000", 
                            "000", "000", "000", "001", "001", "001", "001", "001", 
                            "001", "001", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "111", "111", 
                            "111", "111", "111", "111", "111", "000", "000", "000", 
                            "000", "000", "000", "001", "001", "001", "001", "001", 
                            "001", "001", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "111", "111", 
                            "111", "111", "111", "111", "111", "000", "000", "000", 
                            "000", "000", "000", "001", "001", "001", "001", "001", 
                            "001", "001", "001", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "111", "111", "111", 
                            "111", "111", "111", "111", "111", "000", "000", "000", 
                            "000", "000", "000", "001", "001", "001", "001", "001", 
                            "001", "001", "001", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "010", "010", "010", "010", "010", "010", "010", "010", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "110", "110", "110", 
                            "110", "110", "110", "110", "110", "111", "111", "111", 
                            "111", "111", "111", "111", "111", "000", "000", "000"); 

begin
	process(A, B)
		variable BA: std_logic_vector(8 downto 0);
	begin
    	BA := B & A;
		q <= LUT(to_integer(unsigned(BA)));
	end process;
end architecture;